-- This file should be updated using the script
package file_paths is
    constant loop_program       : string := "/ERROR - RUN THE SCRIPT TO REGENERATED FILE";
    constant calculator_program : string := "/ERROR - RUN THE SCRIPT TO REGENERATED FILE";
    constant max_program        : string := "/ERROR - RUN THE SCRIPT TO REGENERATED FILE";
    constant biglari_program    : string := "/ERROR - RUN THE SCRIPT TO REGENERATED FILE";
end package;