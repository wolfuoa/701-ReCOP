ENTITY flip_flop IS
    PORT MAP(

    );
END ENTITY flip_flop;

ARCHITECTURE arch OF flip_flop IS

    SIGNAL

BEGIN

END arch; -- arch